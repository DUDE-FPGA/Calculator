--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:56:09 04/25/2014
-- Design Name:   
-- Module Name:   C:/Users/James Donnellan/Documents/GitHub/Calculator/fp32_2_bcd/fp32_2_bcdmk2/fp32bcdtest2.vhd
-- Project Name:  fp32_2_bcdmk2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: fp32bcd2
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY fp32bcdtest2 IS
END fp32bcdtest2;
 
ARCHITECTURE behavior OF fp32bcdtest2 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT fp32bcd2
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         start_conv : IN  std_logic;
         ready : OUT  std_logic;
         done_tick : OUT  std_logic;
         fp32 : IN  std_logic_vector(31 downto 0);
         bcds : OUT  std_logic_vector(39 downto 0);
         sign : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal start_conv : std_logic := '0';
   signal fp32 : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal ready : std_logic;
   signal done_tick : std_logic;
   signal bcds : std_logic_vector(39 downto 0);
   signal sign : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: fp32bcd2 PORT MAP (
          clk => clk,
          reset => reset,
          start_conv => start_conv,
          ready => ready,
          done_tick => done_tick,
          fp32 => fp32,
          bcds => bcds,
          sign => sign
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
